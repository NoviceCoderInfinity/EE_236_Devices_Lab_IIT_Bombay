Diode based bridge rectifier

.model diode d()
r1 1 3 1k
d1 1 0 diode
d2 1 2 diode
d3 2 3 diode
d4 0 3 diode

vin 2 0 sin(0 12v 0.05k 0 0)
.tran 0.02ms 40ms
.control
run
plot v(3,1) v(2)
.endc
.end
