Shunt Clipper DC Analysis
r1 1 2 1k
* Defining the diode to be used as the default one
.model diode d()
* Specifying a default diode p n
d1 2 3 diode
*Independent DC Source of 2V
vdc 0 3 dc 2
*Independent DC Source whose voltage is to be varied
vsin 1 0 sin(0 5 1k 0 0)
* Transient analysis
.control
tran 0.02m 10m
set hcopydevtype=postscript
hardcopy Exercise_1_b.ps v(2) v(1)
.endc
.end
