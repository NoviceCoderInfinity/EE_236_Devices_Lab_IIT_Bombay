IV characteristics of Solar Cell

.subckt solar_cell PX NX
*IL is photo generated current (keep only 1 of the next 3 lines, whichever is necessary)
*IL NX TMP dc 0e-3
*IL NX TMP dc 8e-3
IL NX TMP dc 10e-3

d1 TMP NX diode
.model diode d (is=(1e-13) n=1)

d2 TMP NX diode2
.model diode2 d (is=(2e-6) n=2)

*rs TMP PX 0
rs TMP PX 10
*rs TMP PX 30

*rsh TMP NX 5e2
rsh TMP NX 1e3
*rsh TMP NX 5e3

.ends solar_cell

Vin 1 0 dc 0

X1 1 2 solar_cell

r1 2 0 100

.dc Vin -2 2 0.01
.temp 55
.control
run
plot -i(vin) vs {v(1)-v(2)}
wrdata char_10_55C.txt -i(vin) {v(1)-v(2)} 

.endc
.end

